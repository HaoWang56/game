
module altpll0 (
	areset_reset,
	inclk0_clk,
	c0_clk);	

	input		areset_reset;
	input		inclk0_clk;
	output		c0_clk;
endmodule
