// altpll0.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module altpll0 (
		input  wire  areset_reset, // areset.reset
		output wire  c0_clk,       //     c0.clk
		input  wire  inclk0_clk    // inclk0.clk
	);

	altpll0_altpll_0 altpll_0 (
		.clk                (inclk0_clk),   //       inclk_interface.clk
		.reset              (areset_reset), // inclk_interface_reset.reset
		.read               (),             //             pll_slave.read
		.write              (),             //                      .write
		.address            (),             //                      .address
		.readdata           (),             //                      .readdata
		.writedata          (),             //                      .writedata
		.c0                 (c0_clk),       //                    c0.clk
		.areset             (),             //        areset_conduit.export
		.scandone           (),             //           (terminated)
		.scandataout        (),             //           (terminated)
		.locked             (),             //           (terminated)
		.phasedone          (),             //           (terminated)
		.phasecounterselect (4'b0000),      //           (terminated)
		.phaseupdown        (1'b0),         //           (terminated)
		.phasestep          (1'b0),         //           (terminated)
		.scanclk            (1'b0),         //           (terminated)
		.scanclkena         (1'b0),         //           (terminated)
		.scandata           (1'b0),         //           (terminated)
		.configupdate       (1'b0)          //           (terminated)
	);

endmodule
